#include <stdio.h>

int main(int argc, char** argv) {
	printf("hello world");
return 0;
}
